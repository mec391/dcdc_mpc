module MPC_INC_COND(
input i_clk,
input i_rst_n,



	);






endmodule